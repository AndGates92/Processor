library ieee;
use ieee.math_real.all;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;

package ddr2_define_pkg is 

	constant DDR2_CLK_PERIOD	: positive := 1;

end package ddr2_define_pkg;
