library ieee;
use ieee.math_real.all;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;

package common_tb_pkg is 

	constant COMMON_CLK_PERIOD	: integer := 10;

end package common_tb_pkg;
